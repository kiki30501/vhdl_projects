
module mypll (
	inclk,
	ena,
	outclk);	

	input		inclk;
	input		ena;
	output		outclk;
endmodule
